module smoke; initial begin $display("Smoke running"); end endmodule
